`timescale 1ns / 1ps
/******************************************************************************************
* iDEA Soft-Core Processor v1.00
* Copyright (C) by HuiYan Cheah 2012 hycheah1@e.ntu.edu.sg
* School of Computer Engineering
* Nanyang Technological University
*
	* This processor is a proof-of-concept of the usability of the DSP48E1 as
	* the execution unit of a general-purpose processor. It is not a full-blown processor.
	*
	* Description:
	* Instruction Memory of size 512 x 32.
	* Block RAM is inferred through behavioural description.
	* Inferred Block RAM mode is No Change to obtain maximum frequency.
	* Internal output register is enabled.
	* Additional output register in fabric to improve path delay.
	*

******************************************************************************************/
`include "defines.v"

module inst_mem (
	input 						clk,
	input [`im_addr_width-1:0] 	addr_i,
	output reg [31:0] 			dout_o
    );

	reg [31:0] 					rom0 [0:`im_depth-1];
	reg [31:0] 					dout_r0, dout_r1;

	always@ (posedge clk) // No change
	begin
		dout_r0 <= rom0[addr_i];
	end
	
	always@ (posedge clk)
	begin
		dout_r1 <= dout_r0;
		dout_o <= dout_r1;
	end

	initial begin
		//------------cond_s_i_opcod_rd____ra____rb____rc____0
		rom0[0  ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; // 0 nop
		rom0[1  ] = 32'b0110_0_1_11010_00000_0000_0000_0011_0010; //1 movb r0, #0x032 // n = 50
		rom0[2  ] = 32'b0110_0_0_11000_00001_11110_00000_00000_0; //2 mov r1, r30
		rom0[3  ] = 32'b0110_0_1_11010_00010_0000_0000_0000_0001; //3 movb r2, #0x001
		rom0[4  ] = 32'b0110_0_0_11000_00011_11110_00000_00000_0; //4 movb r3, r30
		rom0[5  ] = 32'b0110_0_0_11000_00100_11110_00000_00000_0; //5 mov r4, r30
		rom0[6  ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //6 nop
		rom0[7  ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //7 nop
		rom0[8  ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //8 nop
		rom0[9  ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //9 nop
		rom0[10 ] = 32'b0110_0_0_10010_000000000000000100001____; //10 b  #0x021
		rom0[11 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //11 nop
		rom0[12 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //12 nop
		rom0[13 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //13 nop
		rom0[14 ] = 32'b0110_0_0_00001_00011_00001_00010_00000_0; //14 add r3, r1, r2
		rom0[15 ] = 32'b0110_0_0_11000_00001_00010_00000_00000_0; //15 mov r1, r2
		rom0[16 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //16 nop
		rom0[17 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //17 nop
		rom0[18 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //18 nop
		rom0[19 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //19 nop
		rom0[20 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //20 nop
		rom0[21 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //21 nop
		rom0[22 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //22 nop
		rom0[23 ] = 32'b0110_0_0_11000_00010_00011_00000_00000_0; //23 mov r2, r3
		rom0[24 ] = 32'b0110_0_1_00001_00100_00100_00000_00000_1; //24 add r4, r4, #0x001
		rom0[25 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //25 nop
		rom0[26 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //26 nop
		rom0[27 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //27 nop
		rom0[28 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //28 nop
		rom0[29 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //29 nop
		rom0[30 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //30 nop
		rom0[31 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //31 nop
		rom0[32 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //32 nop
		rom0[33 ] = 32'b0011_1_0_10001_00100_00000_00000001110__; //33 cblt r4, r0, #0x00e (branch target here!)
		rom0[34 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //34 nop
		rom0[35 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //35 nop
		rom0[36 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //36 nop
		rom0[37 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //37 nop
		rom0[38 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //38 nop
		rom0[39 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //39 nop
		rom0[40 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //40 nop
		rom0[41 ] = 32'b0000_0_0_00000_00000_00000_00000_00000_0; //41 nop
		rom0[42	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[43	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[44	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[45	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[46	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[47	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[48	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[49	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[50	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[51	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[52	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[53	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[54	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[55	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[56	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[57	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[58	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[59	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[60	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[61	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[62	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[63	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[64	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[65	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[66	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[67	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[68	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[69	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[70	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[71	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[72	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[73	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[74	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[75	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[76	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[77	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[80	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[81	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[82	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[83	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[84	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[85	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[86	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[87	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[88	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[89	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[90	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[91	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[92	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[93	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[94	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[95	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[96	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[97	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[98	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[99	] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[100] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[101] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[102] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[103] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[104] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[105] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[106] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[107] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[108] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[109] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[110] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[111] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[112] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[113] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[114] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[115] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[116] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[117] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[118] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[119] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[120] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[121] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[122] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[123] =	 32'b0000_0_0_00000_00000_00000_00000_00000_0; //
		rom0[124] = 32'h00000000; rom0[125] = 32'h00000000; rom0[126] = 32'h00000000; rom0[127] = 32'h00000000;
		rom0[128] = 32'h00000000; rom0[129] = 32'h00000000; rom0[130] = 32'h00000000; rom0[131] = 32'h00000000;
		rom0[132] = 32'h00000000; rom0[133] = 32'h00000000; rom0[134] = 32'h00000000; rom0[135] = 32'h00000000;
		rom0[136] = 32'h00000000; rom0[137] = 32'h00000000; rom0[138] = 32'h00000000; rom0[139] = 32'h00000000;
		rom0[140] = 32'h00000000; rom0[141] = 32'h00000000; rom0[142] = 32'h00000000; rom0[143] = 32'h00000000;
		rom0[144] = 32'h00000000; rom0[145] = 32'h00000000; rom0[146] = 32'h00000000; rom0[147] = 32'h00000000;
		rom0[148] = 32'h00000000; rom0[149] = 32'h00000000; rom0[150] = 32'h00000000; rom0[151] = 32'h00000000;
		rom0[152] = 32'h00000000; rom0[153] = 32'h00000000; rom0[154] = 32'h00000000; rom0[155] = 32'h00000000;
		rom0[156] = 32'h00000000; rom0[157] = 32'h00000000; rom0[158] = 32'h00000000; rom0[159] = 32'h00000000;
		rom0[160] = 32'h00000000; rom0[161] = 32'h00000000; rom0[162] = 32'h00000000; rom0[163] = 32'h00000000;
		rom0[164] = 32'h00000000; rom0[165] = 32'h00000000; rom0[166] = 32'h00000000; rom0[167] = 32'h00000000;
		rom0[168] = 32'h00000000; rom0[169] = 32'h00000000; rom0[170] = 32'h00000000; rom0[171] = 32'h00000000;
		rom0[172] = 32'h00000000; rom0[173] = 32'h00000000; rom0[174] = 32'h00000000; rom0[175] = 32'h00000000;
		rom0[176] = 32'h00000000; rom0[177] = 32'h00000000; rom0[178] = 32'h00000000; rom0[179] = 32'h00000000;
		rom0[180] = 32'h00000000; rom0[181] = 32'h00000000; rom0[182] = 32'h00000000; rom0[183] = 32'h00000000;
		rom0[184] = 32'h00000000; rom0[185] = 32'h00000000; rom0[186] = 32'h00000000; rom0[187] = 32'h00000000;
		rom0[188] = 32'h00000000; rom0[189] = 32'h00000000; rom0[190] = 32'h00000000; rom0[191] = 32'h00000000;
		rom0[192] = 32'h00000000; rom0[193] = 32'h00000000; rom0[194] = 32'h00000000; rom0[195] = 32'h00000000;
		rom0[196] = 32'h00000000; rom0[197] = 32'h00000000; rom0[198] = 32'h00000000; rom0[199] = 32'h00000000;
		rom0[200] = 32'h00000000; rom0[201] = 32'h00000000; rom0[202] = 32'h00000000; rom0[203] = 32'h00000000;
		rom0[204] = 32'h00000000; rom0[205] = 32'h00000000; rom0[206] = 32'h00000000; rom0[207] = 32'h00000000;
		rom0[208] = 32'h00000000; rom0[209] = 32'h00000000; rom0[210] = 32'h00000000; rom0[211] = 32'h00000000;
		rom0[212] = 32'h00000000; rom0[213] = 32'h00000000; rom0[214] = 32'h00000000; rom0[215] = 32'h00000000;
		rom0[216] = 32'h00000000; rom0[217] = 32'h00000000; rom0[218] = 32'h00000000; rom0[219] = 32'h00000000;
		rom0[220] = 32'h00000000; rom0[221] = 32'h00000000; rom0[222] = 32'h00000000; rom0[223] = 32'h00000000;
		rom0[224] = 32'h00000000; rom0[225] = 32'h00000000; rom0[226] = 32'h00000000; rom0[227] = 32'h00000000;
		rom0[228] = 32'h00000000; rom0[229] = 32'h00000000; rom0[230] = 32'h00000000; rom0[231] = 32'h00000000;
		rom0[232] = 32'h00000000; rom0[233] = 32'h00000000; rom0[234] = 32'h00000000; rom0[235] = 32'h00000000;
		rom0[236] = 32'h00000000; rom0[237] = 32'h00000000; rom0[238] = 32'h00000000; rom0[239] = 32'h00000000;
		rom0[240] = 32'h00000000; rom0[241] = 32'h00000000; rom0[242] = 32'h00000000; rom0[243] = 32'h00000000;
		rom0[244] = 32'h00000000; rom0[245] = 32'h00000000; rom0[246] = 32'h00000000; rom0[247] = 32'h00000000;
		rom0[248] = 32'h00000000; rom0[249] = 32'h00000000; rom0[250] = 32'h00000000; rom0[251] = 32'h00000000;
		rom0[252] = 32'h00000000; rom0[253] = 32'h00000000; rom0[254] = 32'h00000000; rom0[255] = 32'h00000000;
		rom0[256] = 32'h00000000; rom0[257] = 32'h00000000; rom0[258] = 32'h00000000; rom0[259] = 32'h00000000;
		rom0[260] = 32'h00000000; rom0[261] = 32'h00000000; rom0[262] = 32'h00000000; rom0[263] = 32'h00000000;
		rom0[264] = 32'h00000000; rom0[265] = 32'h00000000; rom0[266] = 32'h00000000; rom0[267] = 32'h00000000;
		rom0[268] = 32'h00000000; rom0[269] = 32'h00000000; rom0[270] = 32'h00000000; rom0[271] = 32'h00000000;
		rom0[272] = 32'h00000000; rom0[273] = 32'h00000000; rom0[274] = 32'h00000000; rom0[275] = 32'h00000000;
		rom0[276] = 32'h00000000; rom0[277] = 32'h00000000; rom0[278] = 32'h00000000; rom0[279] = 32'h00000000;
		rom0[280] = 32'h00000000; rom0[281] = 32'h00000000; rom0[282] = 32'h00000000; rom0[283] = 32'h00000000;
		rom0[284] = 32'h00000000; rom0[285] = 32'h00000000; rom0[286] = 32'h00000000; rom0[287] = 32'h00000000;
		rom0[288] = 32'h00000000; rom0[289] = 32'h00000000; rom0[290] = 32'h00000000; rom0[291] = 32'h00000000;
		rom0[292] = 32'h00000000; rom0[293] = 32'h00000000; rom0[294] = 32'h00000000; rom0[295] = 32'h00000000;
		rom0[296] = 32'h00000000; rom0[297] = 32'h00000000; rom0[298] = 32'h00000000; rom0[299] = 32'h00000000;
		rom0[300] = 32'h00000000; rom0[301] = 32'h00000000; rom0[302] = 32'h00000000; rom0[303] = 32'h00000000;
		rom0[304] = 32'h00000000; rom0[205] = 32'h00000000; rom0[306] = 32'h00000000; rom0[307] = 32'h00000000;
		rom0[308] = 32'h00000000; rom0[309] = 32'h00000000; rom0[310] = 32'h00000000; rom0[311] = 32'h00000000;
		rom0[312] = 32'h00000000; rom0[313] = 32'h00000000; rom0[314] = 32'h00000000; rom0[315] = 32'h00000000;
		rom0[316] = 32'h00000000; rom0[317] = 32'h00000000; rom0[318] = 32'h00000000; rom0[319] = 32'h00000000;
		rom0[320] = 32'h00000000; rom0[321] = 32'h00000000; rom0[322] = 32'h00000000; rom0[323] = 32'h00000000;
		rom0[324] = 32'h00000000; rom0[325] = 32'h00000000; rom0[326] = 32'h00000000; rom0[327] = 32'h00000000;
		rom0[328] = 32'h00000000; rom0[329] = 32'h00000000; rom0[330] = 32'h00000000; rom0[331] = 32'h00000000;
		rom0[332] = 32'h00000000; rom0[333] = 32'h00000000; rom0[334] = 32'h00000000; rom0[335] = 32'h00000000;
		rom0[336] = 32'h00000000; rom0[337] = 32'h00000000; rom0[338] = 32'h00000000; rom0[339] = 32'h00000000;
		rom0[340] = 32'h00000000; rom0[341] = 32'h00000000; rom0[342] = 32'h00000000; rom0[343] = 32'h00000000;
		rom0[344] = 32'h00000000; rom0[345] = 32'h00000000; rom0[346] = 32'h00000000; rom0[347] = 32'h00000000;
		rom0[348] = 32'h00000000; rom0[349] = 32'h00000000; rom0[350] = 32'h00000000; rom0[351] = 32'h00000000;
		rom0[352] = 32'h00000000; rom0[353] = 32'h00000000; rom0[354] = 32'h00000000; rom0[355] = 32'h00000000;
		rom0[356] = 32'h00000000; rom0[357] = 32'h00000000; rom0[358] = 32'h00000000; rom0[359] = 32'h00000000;
		rom0[360] = 32'h00000000; rom0[361] = 32'h00000000; rom0[362] = 32'h00000000; rom0[363] = 32'h00000000;
		rom0[364] = 32'h00000000; rom0[365] = 32'h00000000; rom0[366] = 32'h00000000; rom0[367] = 32'h00000000;
		rom0[368] = 32'h00000000; rom0[369] = 32'h00000000; rom0[370] = 32'h00000000; rom0[371] = 32'h00000000;
		rom0[372] = 32'h00000000; rom0[373] = 32'h00000000; rom0[374] = 32'h00000000; rom0[375] = 32'h00000000;
		rom0[376] = 32'h00000000; rom0[377] = 32'h00000000; rom0[378] = 32'h00000000; rom0[379] = 32'h00000000;
		rom0[380] = 32'h00000000; rom0[381] = 32'h00000000; rom0[382] = 32'h00000000; rom0[383] = 32'h00000000;
		rom0[384] = 32'h00000000; rom0[385] = 32'h00000000; rom0[386] = 32'h00000000; rom0[387] = 32'h00000000;
		rom0[388] = 32'h00000000; rom0[389] = 32'h00000000; rom0[390] = 32'h00000000; rom0[391] = 32'h00000000;
		rom0[392] = 32'h00000000; rom0[393] = 32'h00000000; rom0[394] = 32'h00000000; rom0[395] = 32'h00000000;
		rom0[396] = 32'h00000000; rom0[397] = 32'h00000000; rom0[398] = 32'h00000000; rom0[399] = 32'h00000000;
		rom0[400] = 32'h00000000; rom0[401] = 32'h00000000; rom0[402] = 32'h00000000; rom0[403] = 32'h00000000;
		rom0[404] = 32'h00000000; rom0[405] = 32'h00000000; rom0[406] = 32'h00000000; rom0[407] = 32'h00000000;
		rom0[408] = 32'h00000000; rom0[409] = 32'h00000000; rom0[410] = 32'h00000000; rom0[411] = 32'h00000000;
		rom0[412] = 32'h00000000; rom0[413] = 32'h00000000; rom0[414] = 32'h00000000; rom0[415] = 32'h00000000;
		rom0[416] = 32'h00000000; rom0[417] = 32'h00000000; rom0[418] = 32'h00000000; rom0[419] = 32'h00000000;
		rom0[420] = 32'h00000000; rom0[421] = 32'h00000000; rom0[422] = 32'h00000000; rom0[423] = 32'h00000000;
		rom0[424] = 32'h00000000; rom0[425] = 32'h00000000; rom0[426] = 32'h00000000; rom0[427] = 32'h00000000;
		rom0[428] = 32'h00000000; rom0[429] = 32'h00000000; rom0[430] = 32'h00000000; rom0[431] = 32'h00000000;
		rom0[432] = 32'h00000000; rom0[433] = 32'h00000000; rom0[434] = 32'h00000000; rom0[435] = 32'h00000000;
		rom0[436] = 32'h00000000; rom0[437] = 32'h00000000; rom0[438] = 32'h00000000; rom0[439] = 32'h00000000;
		rom0[440] = 32'h00000000; rom0[441] = 32'h00000000; rom0[442] = 32'h00000000; rom0[443] = 32'h00000000;
		rom0[444] = 32'h00000000; rom0[445] = 32'h00000000; rom0[446] = 32'h00000000; rom0[447] = 32'h00000000;
		rom0[448] = 32'h00000000; rom0[449] = 32'h00000000; rom0[450] = 32'h00000000; rom0[451] = 32'h00000000;
		rom0[452] = 32'h00000000; rom0[453] = 32'h00000000; rom0[454] = 32'h00000000; rom0[455] = 32'h00000000;
		rom0[456] = 32'h00000000; rom0[457] = 32'h00000000; rom0[458] = 32'h00000000; rom0[459] = 32'h00000000;
		rom0[460] = 32'h00000000; rom0[461] = 32'h00000000; rom0[462] = 32'h00000000; rom0[463] = 32'h00000000;
		rom0[464] = 32'h00000000; rom0[465] = 32'h00000000; rom0[466] = 32'h00000000; rom0[467] = 32'h00000000;
		rom0[468] = 32'h00000000; rom0[469] = 32'h00000000; rom0[470] = 32'h00000000; rom0[471] = 32'h00000000;
		rom0[472] = 32'h00000000; rom0[473] = 32'h00000000; rom0[474] = 32'h00000000; rom0[475] = 32'h00000000;
		rom0[476] = 32'h00000000; rom0[477] = 32'h00000000; rom0[478] = 32'h00000000; rom0[479] = 32'h00000000;
		rom0[480] = 32'h00000000; rom0[481] = 32'h00000000; rom0[482] = 32'h00000000; rom0[483] = 32'h00000000;
		rom0[484] = 32'h00000000; rom0[485] = 32'h00000000; rom0[486] = 32'h00000000; rom0[487] = 32'h00000000;
		rom0[488] = 32'h00000000; rom0[489] = 32'h00000000; rom0[490] = 32'h00000000; rom0[491] = 32'h00000000;
		rom0[492] = 32'h00000000; rom0[493] = 32'h00000000; rom0[494] = 32'h00000000; rom0[495] = 32'h00000000;
		rom0[496] = 32'h00000000; rom0[497] = 32'h00000000; rom0[498] = 32'h00000000; rom0[499] = 32'h00000000;
		rom0[500] = 32'h00000000; rom0[501] = 32'h00000000; rom0[502] = 32'h00000000; rom0[503] = 32'h00000000;
		rom0[504] = 32'h00000000; rom0[505] = 32'h00000000; rom0[506] = 32'h00000000; rom0[507] = 32'h00000000;
		rom0[508] = 32'h00000000; rom0[509] = 32'h00000000; rom0[510] = 32'h00000000; rom0[511] = 32'h00000000;
	end

endmodule
